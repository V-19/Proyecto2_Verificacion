`include "ram_dp_ar_aw.v"
`include "sync_fifo.v"
`include "top_hdl.sv"
