// Code your testbench here
// or browse Examples
//`include "tb_core.sv"
`include "tb_top.sv"