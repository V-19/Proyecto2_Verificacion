// Code your design here
`include "sdrc_bank_ctl.v"
`include "sdrc_bank_fsm.v"
`include "sdrc_bs_convert.v"
`include "sdrc_core.v"
`include "sdrc_req_gen.v"
`include "sdrc_top.v"
`include "sdrc_xfr_ctl.v"
`include "sdrc_define.v"
`include "async_fifo.v"
`include "sync_fifo.v"
`include "wb2sdrc.v"
`include "mt48lc2m32b2.v"
//`include "IS42VM16400K.V"
`include "mt48lc8m8a2.v"
`include "top_hdl.sv"